`include "datapath.vh"

module skintone_datapath
(
	input				clk, 
	input 				rst,
	input 	[23:0]			pixel_datain, 
	input				pixel_datain_valid,
	input				pixel_datain_ready,
	output	[7:0]			result_dataout,
	output				result_dataout_valid,
	output				result_dataout_ready
);



endmodule