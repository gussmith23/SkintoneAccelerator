module transcx
(
	input 		clk,
	input 	[7:0]	Cx,
	input 	[7:0]	Y,
	output	[7:0]	transcx
);

endmodule;