`include "datapath.h"

module fp_mult
(

)